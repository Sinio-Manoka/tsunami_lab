netcdf 03_tsunami_lab { // example showing how output of the tsunami lab might look like
dimensions:
    x = 3;
    y = 8;
    time = unlimited;
variables:
    float x(x);
      x:units = "meters";
      x:axis = "X";
    float y(y);
      x:units = "meters";
      x:axis = "Y";
    float time(time);
      time:units = "seconds";
    float b(y, x);
      b:units = "meters";
    float h(time, y, x);
      h:units = "meters";
    // TODO: hu and hv go here
// global attributes
    :title = "Example output of the tsunami lab's solver";
    :summary = "Example output for the solvers of the tsunami lab at Friedrich Schiller University Jena. Further information is available from: https://scalable.uni-jena.de";
data:
  x = 1.5, 2.0, 2.5;
  y = 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0;
  time = 0.0, 25.0, 50.0;
  b =  -2,  -3,  -5,
       -7, -11, -13,
      -17, -19, -23,
      -29, -31, -37,
      -41, -43, -47,
      -53, -59, -61,
      -67, -71, -73,
      -79, -83, -89;
  h =  2,  3,  5,
       7, 11, 13,
      17, 19, 23,
      29, 31, 37,
      41, 43, 47,
      53, 59, 61,
      67, 71, 73,
      79, 83, 89,

       2,    3,    5,
       7,   11,   13,
      17,   19,   23,
      29,   31,   37,
      41.5, 43.5, 47.5,
      53.5, 60,   61.5,
      67.5, 71.5, 73.5,
      79,   83,   89,

       2,     3,     5,
       7,    11,    13,
      17,    19,    23,
      29.05, 31.1,  37.05,
      41.25, 43.25, 47.25,
      53.25, 60.5,  61.25,
      67.25, 71.25, 73.25,
      79.05, 83.1,  89.05;
}